/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Module: RL_LJ_Intergrated_Top.v
//
//	Function:
//				Integrated top module holding all the cells in the simulation space
//
//	Purpose:
//				For real simulation with all the dataset
//				Timing testing with the integrated system
//
// Data Organization:
//				Address 0 for each cell module: # of particles in the cell.
//				MSB-LSB: {posz, posy, posx}
//
// Used by:
//				NA
//
// Dependency:
//				RL_LJ_Evaluation_Unit.v
//				Particle_Pair_Gen_HalfShell.v
//				Motion_Update.v
//				cell_x_y_z.v
//				Force_Cache_x_y_z.v
//				Velocity_Cache_x_y_z.v
//
// Testbench:
//				TBD
//
// Timing:
//				TBD
//
// Created by:
//				Chen Yang's Script (Gen_Sim_Top.cpp)
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module RL_LJ_Intergrated_Top
#(
	parameter DATA_WIDTH 					= 32,
	// Simulation parameters
	parameter TIME_STEP 						= 32'h27101D7D,							// 2fs time step
	// The home cell this unit is working on
	parameter CELL_X							= 4'd2,
	parameter CELL_Y							= 4'd2,
	parameter CELL_Z							= 4'd2,
	// High level parameters
	parameter NUM_EVAL_UNIT					= 1,									// # of evaluation units in the design
	// Dataset defined parameters	parameter MAX_CELL_COUNT_PER_DIM 		= 5,									// Maximum cell count among the 3 dimensions
	parameter NUM_NEIGHBOR_CELLS				= 13,									// # of neighbor cells per home cell, for Half-shell method, is 13
	parameter CELL_ID_WIDTH					= 3,									// log(NUM_NEIGHBOR_CELLS)
	parameter MAX_CELL_PARTICLE_NUM			= 290,									// The maximum # of particles can be in a cell
	parameter CELL_ADDR_WIDTH				= 9,									// log(MAX_CELL_PARTICLE_NUM)
	parameter PARTICLE_ID_WIDTH				= CELL_ID_WIDTH*3+CELL_ADDR_WIDTH,		// # of bit used to represent particle ID, 9*9*7 cells, each 4-bit, each cell have max of 220 particles, 8-bit
	// Filter parameters	parameter NUM_FILTER						= 8,		//4
	parameter ARBITER_MSB 					= 128,	//8								// 2^(NUM_FILTER-1)
	parameter FILTER_BUFFER_DEPTH 			= 32,
	parameter FILTER_BUFFER_ADDR_WIDTH		= 5,
	parameter CUTOFF_2 						= 32'h43100000,							// (12^2=144 in IEEE floating point)
	// Force Evaluation parameters	parameter SEGMENT_NUM					= 14,
	parameter SEGMENT_WIDTH					= 4,
	parameter BIN_NUM						= 256,
	parameter BIN_WIDTH						= 8,
	parameter LOOKUP_NUM						= SEGMENT_NUM * BIN_NUM,				// SEGMENT_NUM * BIN_NUM
	parameter LOOKUP_ADDR_WIDTH				= SEGMENT_WIDTH + BIN_WIDTH,			// log LOOKUP_NUM / log 2
	// Force (accmulation) cache parameters	parameter FORCE_CACHE_BUFFER_DEPTH		= 16,									// Force cache input buffer depth, for partial force accumulation
	parameter FORCE_CACHE_BUFFER_ADDR_WIDTH	= 4										// log(FORCE_CACHE_BUFFER_DEPTH) / log 2
)
(
	input clk,
	input rst,
	input start,
	// These are all temp output ports	output [NUM_EVAL_UNIT*PARTICLE_ID_WIDTH-1:0] ref_particle_id,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] ref_LJ_Force_X,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] ref_LJ_Force_Y,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] ref_LJ_Force_Z,
	output [NUM_EVAL_UNIT-1:0] ref_forceoutput_valid,
	output [NUM_EVAL_UNIT*PARTICLE_ID_WIDTH-1:0] neighbor_particle_id,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] neighbor_LJ_Force_X,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] neighbor_LJ_Force_Y,
	output [NUM_EVAL_UNIT*DATA_WIDTH-1:0] neighbor_LJ_Force_Z,
	output [NUM_EVAL_UNIT-1:0] neighbor_forceoutput_valid,
	// Done signals
	// When entire home cell is done processing, this will keep high until the next time 'start' signal turn high
	output out_home_cell_evaluation_done,
	// When motion update is done processing, remain high until the next motion update starts
	output out_motion_update_done,
	// Dummy signal selecting which cell is the home cell
	// Need a logic to replace this, generate by out_Motion_Update_cur_cell
	input [3:0] in_sel,
	// Dummy output for motion update
	output [3*CELL_ID_WIDTH-1:0] out_Motion_Update_cur_cell
);

	Pos_Cache_1_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(1),
		.CELL_X(1),
	)
	cell_1_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(1),
		.CELL_X(2),
	)
	cell_1_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(1),
		.CELL_X(3),
	)
	cell_1_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(1),
		.CELL_X(4),
	)
	cell_1_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_1_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(1),
		.CELL_X(5),
	)
	cell_1_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(2),
		.CELL_X(1),
	)
	cell_1_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(2),
		.CELL_X(2),
	)
	cell_1_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(2),
		.CELL_X(3),
	)
	cell_1_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(2),
		.CELL_X(4),
	)
	cell_1_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_2_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(2),
		.CELL_X(5),
	)
	cell_1_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(3),
		.CELL_X(1),
	)
	cell_1_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(3),
		.CELL_X(2),
	)
	cell_1_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(3),
		.CELL_X(3),
	)
	cell_1_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(3),
		.CELL_X(4),
	)
	cell_1_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_3_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(3),
		.CELL_X(5),
	)
	cell_1_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(4),
		.CELL_X(1),
	)
	cell_1_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(4),
		.CELL_X(2),
	)
	cell_1_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(4),
		.CELL_X(3),
	)
	cell_1_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(4),
		.CELL_X(4),
	)
	cell_1_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_4_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(4),
		.CELL_X(5),
	)
	cell_1_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_5_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(5),
		.CELL_X(1),
	)
	cell_1_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_5_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(5),
		.CELL_X(2),
	)
	cell_1_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_5_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(5),
		.CELL_X(3),
	)
	cell_1_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_5_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(5),
		.CELL_X(4),
	)
	cell_1_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_1_5_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_X(5),
		.CELL_X(5),
	)
	cell_1_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(1),
		.CELL_X(1),
	)
	cell_2_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(1),
		.CELL_X(2),
	)
	cell_2_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(1),
		.CELL_X(3),
	)
	cell_2_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(1),
		.CELL_X(4),
	)
	cell_2_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_1_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(1),
		.CELL_X(5),
	)
	cell_2_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(2),
		.CELL_X(1),
	)
	cell_2_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(2),
		.CELL_X(2),
	)
	cell_2_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(2),
		.CELL_X(3),
	)
	cell_2_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(2),
		.CELL_X(4),
	)
	cell_2_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_2_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(2),
		.CELL_X(5),
	)
	cell_2_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(3),
		.CELL_X(1),
	)
	cell_2_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(3),
		.CELL_X(2),
	)
	cell_2_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(3),
		.CELL_X(3),
	)
	cell_2_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(3),
		.CELL_X(4),
	)
	cell_2_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_3_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(3),
		.CELL_X(5),
	)
	cell_2_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(4),
		.CELL_X(1),
	)
	cell_2_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(4),
		.CELL_X(2),
	)
	cell_2_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(4),
		.CELL_X(3),
	)
	cell_2_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(4),
		.CELL_X(4),
	)
	cell_2_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_4_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(4),
		.CELL_X(5),
	)
	cell_2_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_5_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(5),
		.CELL_X(1),
	)
	cell_2_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_5_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(5),
		.CELL_X(2),
	)
	cell_2_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_5_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(5),
		.CELL_X(3),
	)
	cell_2_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_5_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(5),
		.CELL_X(4),
	)
	cell_2_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_2_5_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_X(5),
		.CELL_X(5),
	)
	cell_2_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(1),
		.CELL_X(1),
	)
	cell_3_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(1),
		.CELL_X(2),
	)
	cell_3_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(1),
		.CELL_X(3),
	)
	cell_3_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(1),
		.CELL_X(4),
	)
	cell_3_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_1_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(1),
		.CELL_X(5),
	)
	cell_3_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(2),
		.CELL_X(1),
	)
	cell_3_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(2),
		.CELL_X(2),
	)
	cell_3_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(2),
		.CELL_X(3),
	)
	cell_3_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(2),
		.CELL_X(4),
	)
	cell_3_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_2_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(2),
		.CELL_X(5),
	)
	cell_3_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(3),
		.CELL_X(1),
	)
	cell_3_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(3),
		.CELL_X(2),
	)
	cell_3_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(3),
		.CELL_X(3),
	)
	cell_3_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(3),
		.CELL_X(4),
	)
	cell_3_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_3_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(3),
		.CELL_X(5),
	)
	cell_3_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(4),
		.CELL_X(1),
	)
	cell_3_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(4),
		.CELL_X(2),
	)
	cell_3_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(4),
		.CELL_X(3),
	)
	cell_3_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(4),
		.CELL_X(4),
	)
	cell_3_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_4_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(4),
		.CELL_X(5),
	)
	cell_3_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_5_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(5),
		.CELL_X(1),
	)
	cell_3_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_5_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(5),
		.CELL_X(2),
	)
	cell_3_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_5_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(5),
		.CELL_X(3),
	)
	cell_3_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_5_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(5),
		.CELL_X(4),
	)
	cell_3_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_3_5_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_X(5),
		.CELL_X(5),
	)
	cell_3_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(1),
		.CELL_X(1),
	)
	cell_4_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(1),
		.CELL_X(2),
	)
	cell_4_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(1),
		.CELL_X(3),
	)
	cell_4_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(1),
		.CELL_X(4),
	)
	cell_4_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_1_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(1),
		.CELL_X(5),
	)
	cell_4_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(2),
		.CELL_X(1),
	)
	cell_4_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(2),
		.CELL_X(2),
	)
	cell_4_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(2),
		.CELL_X(3),
	)
	cell_4_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(2),
		.CELL_X(4),
	)
	cell_4_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_2_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(2),
		.CELL_X(5),
	)
	cell_4_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(3),
		.CELL_X(1),
	)
	cell_4_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(3),
		.CELL_X(2),
	)
	cell_4_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(3),
		.CELL_X(3),
	)
	cell_4_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(3),
		.CELL_X(4),
	)
	cell_4_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_3_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(3),
		.CELL_X(5),
	)
	cell_4_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(4),
		.CELL_X(1),
	)
	cell_4_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(4),
		.CELL_X(2),
	)
	cell_4_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(4),
		.CELL_X(3),
	)
	cell_4_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(4),
		.CELL_X(4),
	)
	cell_4_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_4_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(4),
		.CELL_X(5),
	)
	cell_4_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_5_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(5),
		.CELL_X(1),
	)
	cell_4_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_5_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(5),
		.CELL_X(2),
	)
	cell_4_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_5_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(5),
		.CELL_X(3),
	)
	cell_4_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_5_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(5),
		.CELL_X(4),
	)
	cell_4_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_4_5_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_X(5),
		.CELL_X(5),
	)
	cell_4_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(1),
		.CELL_X(1),
	)
	cell_5_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(1),
		.CELL_X(2),
	)
	cell_5_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(1),
		.CELL_X(3),
	)
	cell_5_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(1),
		.CELL_X(4),
	)
	cell_5_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_1_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(1),
		.CELL_X(5),
	)
	cell_5_1_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(2),
		.CELL_X(1),
	)
	cell_5_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(2),
		.CELL_X(2),
	)
	cell_5_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(2),
		.CELL_X(3),
	)
	cell_5_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(2),
		.CELL_X(4),
	)
	cell_5_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_2_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(2),
		.CELL_X(5),
	)
	cell_5_2_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(3),
		.CELL_X(1),
	)
	cell_5_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(3),
		.CELL_X(2),
	)
	cell_5_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(3),
		.CELL_X(3),
	)
	cell_5_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(3),
		.CELL_X(4),
	)
	cell_5_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_3_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(3),
		.CELL_X(5),
	)
	cell_5_3_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(4),
		.CELL_X(1),
	)
	cell_5_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(4),
		.CELL_X(2),
	)
	cell_5_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(4),
		.CELL_X(3),
	)
	cell_5_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(4),
		.CELL_X(4),
	)
	cell_5_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_4_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(4),
		.CELL_X(5),
	)
	cell_5_4_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_5_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(5),
		.CELL_X(1),
	)
	cell_5_5_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_5_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(5),
		.CELL_X(2),
	)
	cell_5_5_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_5_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(5),
		.CELL_X(3),
	)
	cell_5_5_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_5_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(5),
		.CELL_X(4),
	)
	cell_5_5_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

	Pos_Cache_5_5_5
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(MAX_CELL_PARTICLE_NUM),
		.ADDR_WIDTH(CELL_ADDR_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(5),
		.CELL_X(5),
		.CELL_X(5),
	)
	cell_5_5_5
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? Motion_Update_position_read_addr : FSM_to_Cell_read_addr[1*CELL_ADDR_WIDTH-1:0*CELL_ADDR_WIDTH]),
		.in_data(Motion_Update_out_position_data),
		.in_data_dst_cell(Motion_Update_dst_cell),					// The destination cell for the incoming data
		.in_data_valid(Motion_Update_out_position_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? Motion_Update_position_read_en : FSM_to_Cell_rden),
		.out_particle_info(Position_Cache_readout_position[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	)

endmodule
